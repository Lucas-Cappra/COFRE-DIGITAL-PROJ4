LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY COMPARADOR IS
    Port(
        A, B : IN STD_LOGIC;
        GT, LT, EQ: OUT STD_LOGIC
    );
END COMPARADOR;

ARCHITECTURE COMPARADOR OF COMPARADOR IS
SIGNAL GT_AUX, LT_AUX: STD_LOGIC;
BEGIN

GT_AUX <= A AND NOT(B);
LT_AUX <= NOT(A) AND B;

GT <= GT_AUX;
LT <= LT_AUX;
EQ <= NOT (GT_AUX OR LT_AUX);

END ARCHITECTURE COMPARADOR;