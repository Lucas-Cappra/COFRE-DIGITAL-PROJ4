LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY COMPARADOR_18BITS IS
    Port(
        A, B: IN STD_LOGIC_VECTOR (17 DOWNTO 0);
        GT, LT, EQ: OUT STD_LOGIC
    );
END COMPARADOR_18BITS;

ARCHITECTURE COMPARADOR_18BITS OF COMPARADOR_18BITS IS

COMPONENT COMPARADOR IS
    Port(
        A, B: IN STD_LOGIC;
        GT, LT, EQ: OUT STD_LOGIC
    );
END COMPONENT COMPARADOR;


SIGNAL GT0, LT0, EQ0, GT1, LT1, EQ1, GT2, LT2, EQ2: STD_LOGIC;
SIGNAL GT3, LT3, EQ3, GT4, LT4, EQ4, GT5, LT5, EQ5: STD_LOGIC;
SIGNAL GT6, LT6, EQ6, GT7, LT7, EQ7, GT8, LT8, EQ8: STD_LOGIC;
SIGNAL GT9, LT9, EQ9, GT10, LT10, EQ10, GT11, LT11, EQ11: STD_LOGIC;
SIGNAL GT12, LT12, EQ12, GT13, LT13, EQ13, GT14, LT14, EQ14: STD_LOGIC;
SIGNAL GT15, LT15, EQ15, GT16, LT16, EQ16, GT17, LT17, EQ17: STD_LOGIC;

SIGNAL GT_AUX: STD_LOGIC;

BEGIN
C0: COMPARADOR PORT MAP (A(0), B(0), GT0, LT0, EQ0);
C1: COMPARADOR PORT MAP (A(1), B(1), GT1, LT1, EQ1);
C2: COMPARADOR PORT MAP (A(2), B(2), GT2, LT2, EQ2);
C3: COMPARADOR PORT MAP (A(3), B(3), GT3, LT3, EQ3);
C4: COMPARADOR PORT MAP (A(4), B(4), GT4, LT4, EQ4);
C5: COMPARADOR PORT MAP (A(5), B(5), GT5, LT5, EQ5);
C6: COMPARADOR PORT MAP (A(6), B(6), GT6, LT6, EQ6);
C7: COMPARADOR PORT MAP (A(7), B(7), GT7, LT7, EQ7);
C8: COMPARADOR PORT MAP (A(8), B(8), GT8, LT8, EQ8);
C9: COMPARADOR PORT MAP (A(9), B(9), GT9, LT9, EQ9);
C10: COMPARADOR PORT MAP(A(10), B(10), GT10, LT10, EQ10);
C11: COMPARADOR PORT MAP(A(11), B(11), GT11, LT11, EQ11);
C12: COMPARADOR PORT MAP(A(12), B(12), GT12, LT12, EQ12);
C13: COMPARADOR PORT MAP(A(13), B(13), GT13, LT13, EQ13);
C14: COMPARADOR PORT MAP(A(14), B(14), GT14, LT14, EQ14);
C15: COMPARADOR PORT MAP(A(15), B(15), GT15, LT15, EQ15);
C16: COMPARADOR PORT MAP(A(16), B(16), GT16, LT16, EQ16);
C17: COMPARADOR PORT MAP(A(17), B(17), GT17, LT17, EQ17);

GT_AUX <= GT0 OR GT1 OR GT2 OR GT3 OR GT4 OR GT5 OR GT6 OR GT7 OR GT8 OR GT9 OR GT10 OR GT11 OR GT12 OR GT13 OR GT14 OR GT15 OR GT16 OR GT17;

GT <= GT_AUX;
LT <= NOT(GT_AUX);
EQ <= (EQ0 AND EQ1 AND EQ2 AND EQ3 AND EQ4 AND EQ5 AND EQ6 AND EQ7 AND EQ8 AND EQ9 AND EQ10 AND EQ11 AND EQ12 AND EQ13 AND EQ14 AND EQ15 AND EQ16 AND EQ17);

END ARCHITECTURE COMPARADOR_18BITS;
