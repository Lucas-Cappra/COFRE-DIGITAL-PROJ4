LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY LED_RGB IS
	PORT(
		PWR, CONTADOR_20, LOAD: IN STD_LOGIC;
		R, G, B: OUT STD_LOGIC
);
END ENTITY LED_RGB;

ARCHITECTURE LEDS OF LED_RGB IS

	SIGNAL G_AUX, B_AUX: STD_LOGIC;

BEGIN

G_AUX <= CONTADOR_20 AND NOT(B_AUX) AND NOT(PWR);
B_AUX <= PWR XOR LOAD;

R <= NOT(PWR) AND NOT(G_AUX) AND NOT(B_AUX);
G <= G_AUX;
B <= B_AUX;

END ARCHITECTURE LEDS;