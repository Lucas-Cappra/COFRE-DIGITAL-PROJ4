LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY MAQUINA_DE_ESTADOS is
    Port(
        PWR, ADD: IN STD_LOGIC;
	CK: IN STD_LOGIC;
	PWD: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	S: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        PWD_COMP: OUT STD_LOGIC
    );
END MAQUINA_DE_ESTADOS;

ARCHITECTURE COFRE OF MAQUINA_DE_ESTADOS IS
	COMPONENT mde_moore1p is
	port (ck, rst, PWR : in  std_logic;
		ADD, TEMP5, TEMP20, PWD_LEN, PWD_CMP: in  std_logic;
        	q : out std_logic_vector(2 downto 0));
	END COMPONENT mde_moore1p;
	
	COMPONENT SENHA IS 
	Port(
        	PWR, ADD: IN STD_LOGIC;
		PWD: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		S: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        	PWD_COMP: OUT STD_LOGIC
	);
	END COMPONENT SENHA;
	
	COMPONENT LED_RGB IS
	PORT(
		PWR, CONTADOR_20, LOAD: IN STD_LOGIC;
		R, G, B: OUT STD_LOGIC
	);
	END COMPONENT LED_RGB;

	COMPONENT CONTADOR_SENHA IS 
	PORT(
		S: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		CK_IN, CLR, SET: IN STD_LOGIC;
		PWD_LEN: OUT STD_LOGIC  	 		
	);
	END COMPONENT CONTADOR_SENHA;

	COMPONENT TEMPORIZADOR is
    	PORT(
        	S: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		CK: IN STD_LOGIC;
        	TEMP5, TEMP20: OUT STD_LOGIC
    	);
	END COMPONENT TEMPORIZADOR;

	COMPONENT ACESSO IS
	PORT(
		S: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		CLK, CLR, SET: IN STD_LOGIC;
		S_OUT: OUT STD_LOGIC
	);
	END COMPONENT ACESSO;
	
	SIGNAL PWD_COMP_AUX, TEMP20_AUX, TEMP5_AUX, PWD_LEN_AUX: STD_LOGIC;
	SIGNAL R_AUX, G_AUX, B_AUX: STD_LOGIC;
	SIGNAL RST : STD_LOGIC;
	SIGNAL S_AUX: STD_LOGIC_VECTOR (2 DOWNTO 0);

BEGIN

MDE: mde_moore1p PORT MAP (CK, RST, PWR, ADD, TEMP5_AUX, TEMP20_AUX, PWD_LEN_AUX, PWD_COMP_AUX,S_AUX);

S <= S_AUX;

REG_SENHA: SENHA PORT MAP (PWR, ADD, PWD, S_AUX, PWD_COMP_AUX);
TEMP: TEMPORIZADOR PORT MAP (S_AUX, CK, TEMP5_AUX, TEMP20_AUX);
CONT_SENHA: CONTADOR_SENHA PORT MAP (S_AUX,CK,'1', '1', PWD_LEN_AUX);
RGB: LED_RBG PORT MAP (PWR, TEMP20_AUX, ADD, R_AUX, G_AUX, B_AUX);
ACC:  ACESSO PORT MAP (S_AUX, CK, '1', '1', S_ACESSO);
  
  



END ARCHITECTURE;
