LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY CONTADOR_SENHA IS 
	PORT(
		S: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		CK_IN, CLR, SET: IN STD_LOGIC;
		PWD_LEN: OUT STD_LOGIC  		
);
END CONTADOR_SENHA;


ARCHITECTURE CONTADOR_SENHA OF CONTADOR_SENHA IS
	COMPONENT ffd is
   		PORT (ck, clr, set, d : in  std_logic;
                       q : out std_logic);
	END COMPONENT ffd;

	COMPONENT Somador_Completo is
		Port(
        	A_SC, B_SC, CI_SC: IN STD_LOGIC;
        	S_SC, CO_SC: OUT STD_LOGIC
    	);
	END COMPONENT  Somador_Completo;

	COMPONENT mux_2x1 is
	Port (
        	A, B : in  STD_LOGIC;
        	C    : in  STD_LOGIC;
        	Y    : out STD_LOGIC
    	);
	END COMPONENT mux_2x1;

	COMPONENT COMPARADOR_3BITS IS
    	Port(
        	A, B: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
        	GT, LT, EQ: OUT STD_LOGIC
    	);
	END COMPONENT COMPARADOR_3BITS;
	
	SIGNAL Q1_AUX, Q2_AUX, FFD_AUX, S1, COUT_1, S2, COUT_2: STD_LOGIC;
	SIGNAL GT, LT, EQ, MUX_AUX: STD_LOGIC;
	SIGNAL S1_AUX, S2_AUX: STD_LOGIC;
	--SIGNAL CK_OUT: STD_LOGIC;

BEGIN

COMP: COMPARADOR_3BITS PORT MAP (S,"100",GT, LT, EQ);

ENABLE: MUX_2X1 PORT MAP ('0', '1', EQ, MUX_AUX);

FFD_1: FFD PORT MAP (CK_IN, CLR, SET, MUX_AUX, Q1_AUX);
FFD_2: FFD PORT MAP (CK_IN, CLR, SET, Q1_AUX, Q2_AUX);

FFD_AUX <= Q1_AUX AND Q2_AUX;


FFD_SOMA1: FFD PORT MAP (CK_IN, CLR, SET, S1, S1_AUX);
FFD_SOMA2: FFD PORT MAP (CK_IN, CLR, SET, S2, S2_AUX);

SS1: SOMADOR_COMPLETO PORT MAP (FFD_AUX, S1_AUX , '0', S1, COUT_1);
SS2: SOMADOR_COMPLETO PORT MAP (S2_AUX,'0', COUT_1, S2, COUT_2);

PWD_LEN <= (S1_AUX AND '1') AND (S2_AUX AND '1');

 END ARCHITECTURE; 
